module afe_configure
       (
         input clk, reset_n,
         input miso,
         output pdn,
         output cs_n,
         output mosi,
         output device_reset,
         output configure_done
       );

endmodule
